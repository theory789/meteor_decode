/home/sammy/shit/lrpt_decoder/hdl/viterbi.sv