/home/sammy/shit/lrpt_decoder/hdl/tbu.sv