/home/sammy/shit/lrpt_decoder/hdl/bmu.sv