/home/sammy/shit/lrpt_decoder/hdl/acs_but.sv